`timescale 1ns / 1ps
module IOBUF#(
    parameter DRIVE = 12,
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW = "SLOW"
)(
    input           I,
    inout           IO,
    output          O,
    input           T
    );

    // NULL MODULE

endmodule